/*******************************************************************************
  Copyright 2019 Benjamin Devlin

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/

module async_mult #(
  parameter BITS
) (
  input [BITS-1:0]          i_dat_a,
  input [BITS-1:0]          i_dat_b,
  output logic [2*BITS-1:0] o_dat
);

always_comb
  o_dat = i_dat_a * i_dat_b;

endmodule