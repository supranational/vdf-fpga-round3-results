/*******************************************************************************
  Copyright 2019 Steve Golson

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/

(* use_dsp = "yes" *)
module mult_26x17 (x,y,p);

   input  [26-1:0]      x;
   input  [17-1:0]      y;
   output [(26+17)-1:0] p;

   assign p = x * y;

endmodule

